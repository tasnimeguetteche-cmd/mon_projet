* Caractérisation de la consommation statique - xor3_1
.title Static Power Characterization xor3_1

* ============================================
* Conditions de fonctionnement (PVT)
* ============================================
* Process: tt (typical-typical)
.lib "~/.ciel/sky130A/libs.tech/ngspice/sky130.lib.spice" tt

* Voltage: 1.8V (nominal)
.param VDD_VAL = 1.8

* Temperature: 25°C (nominal)
.temp 25

* ============================================
* Inclusion des cellules standard
* ============================================
.include "~/.ciel/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

* ============================================
* Alimentations globales
* ============================================
.global VPWR VGND VNB VPB
VVPWR VPWR 0 DC {VDD_VAL}
VVGND VGND 0 DC 0
VVNB VNB 0 DC 0
VVPB VPB 0 DC {VDD_VAL}

* ============================================
* Instance de la cellule XOR3_1
* ============================================
X1 A B C VGND VNB VPB VPWR Y sky130_fd_sc_hd__xor3_1

* ============================================
* Stimuli des entrées - Séquence des 8 états
* Transition lente entre les états pour stabilisation
* ============================================
VA A VGND PWL(
+ 0n     0
+ 10n    0
+ 11n    0
+ 20n    0
+ 21n    0
+ 30n    0
+ 31n    0
+ 40n    0
+ 41n    1.8
+ 50n    1.8
+ 51n    1.8
+ 60n    1.8
+ 61n    1.8
+ 70n    1.8
+ 71n    1.8
+ 80n    1.8
+ )

VB B VGND PWL(
+ 0n     0
+ 10n    0
+ 11n    0
+ 20n    0
+ 21n    1.8
+ 30n    1.8
+ 31n    1.8
+ 40n    1.8
+ 41n    0
+ 50n    0
+ 51n    0
+ 60n    0
+ 61n    1.8
+ 70n    1.8
+ 71n    1.8
+ 80n    1.8
+ )

VC C VGND PWL(
+ 0n     0
+ 10n    0
+ 11n    1.8
+ 20n    1.8
+ 21n    0
+ 30n    0
+ 31n    1.8
+ 40n    1.8
+ 41n    0
+ 50n    0
+ 51n    1.8
+ 60n    1.8
+ 61n    0
+ 70n    0
+ 71n    1.8
+ 80n    1.8
+ )

* ============================================
* Options de simulation
* ============================================
.option POST
.option NOMOD

* ============================================
* Analyse transitoire pour passer par tous les états
* ============================================
.tran 0.1n 85n

* ============================================
* Mesures de la consommation statique pour chaque état
* Mesure au milieu de chaque état stable (à t=5n de chaque début)
* ============================================

* État 000 (A=0, B=0, C=0) -> Y=0
.measure tran I_static_000 FIND I(VVPWR) AT=5n
.measure tran P_static_000 PARAM='abs(I_static_000)*VDD_VAL'

* État 001 (A=0, B=0, C=1) -> Y=1
.measure tran I_static_001 FIND I(VVPWR) AT=15n
.measure tran P_static_001 PARAM='abs(I_static_001)*VDD_VAL'

* État 010 (A=0, B=1, C=0) -> Y=1
.measure tran I_static_010 FIND I(VVPWR) AT=25n
.measure tran P_static_010 PARAM='abs(I_static_010)*VDD_VAL'

* État 011 (A=0, B=1, C=1) -> Y=0
.measure tran I_static_011 FIND I(VVPWR) AT=35n
.measure tran P_static_011 PARAM='abs(I_static_011)*VDD_VAL'

* État 100 (A=1, B=0, C=0) -> Y=1
.measure tran I_static_100 FIND I(VVPWR) AT=45n
.measure tran P_static_100 PARAM='abs(I_static_100)*VDD_VAL'

* État 101 (A=1, B=0, C=1) -> Y=0
.measure tran I_static_101 FIND I(VVPWR) AT=55n
.measure tran P_static_101 PARAM='abs(I_static_101)*VDD_VAL'

* État 110 (A=1, B=1, C=0) -> Y=0
.measure tran I_static_110 FIND I(VVPWR) AT=65n
.measure tran P_static_110 PARAM='abs(I_static_110)*VDD_VAL'

* État 111 (A=1, B=1, C=1) -> Y=1
.measure tran I_static_111 FIND I(VVPWR) AT=75n
.measure tran P_static_111 PARAM='abs(I_static_111)*VDD_VAL'

* ============================================
* Calcul de la consommation statique moyenne
* ============================================
.measure tran P_static_avg PARAM='(P_static_000+P_static_001+P_static_010+P_static_011+P_static_100+P_static_101+P_static_110+P_static_111)/8'

* ============================================
* Commandes de contrôle
* ============================================
.control
run

* Affichage des signaux
plot V(A)+6 V(B)+4 V(C)+2 V(Y) title 'Static Power - Input States'
plot I(VVPWR)*1e9 title 'Leakage Current (nA)'

* Affichage des résultats
echo "=========================================="
echo "STATIC POWER CHARACTERIZATION - XOR3_1"
echo "=========================================="
echo "Process: tt | Voltage: 1.8V | Temperature: 25°C"
echo "=========================================="
print P_static_000 P_static_001 P_static_010 P_static_011
print P_static_100 P_static_101 P_static_110 P_static_111
echo "=========================================="
print P_static_avg
echo "=========================================="

* Sauvegarde
write static_xor3_1.raw

.endc

.end
