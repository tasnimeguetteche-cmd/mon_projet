.param VDD=1.8
.param L=1.5e-07
.param W_N=2.3599999999999977e-06
.param W_P=3.981663219440153e-06
