* Test Porte ET 
.title Porte ET

.include "params.spice"

.param VDD_VAL = 1.8

* ============================================
* Alimentations
* ============================================
VVDD vdd 0 DC {VDD_VAL}

* ============================================
* PORTE ET CMOS (NAND + INV)
* ============================================
.model nfet_simple nmos (level=54 version=4.5)
.model pfet_simple pmos (level=54 version=4.5)

* --- Étage NAND ---
* On relie A et B ensemble au signal "in" pour le test
MN0 n_nand in node_int 0 nfet_simple W={W_N} L={L}
MN1 node_int in 0 0       nfet_simple W={W_N} L={L}

MP0 n_nand in vdd vdd     pfet_simple W={W_P} L={L}
MP1 n_nand in vdd vdd     pfet_simple W={W_P} L={L}

* --- Étage INVERSEUR ---
* La sortie finale est "out" pour correspondre à vos mesures
MNinv out n_nand 0 0        nfet_simple W={W_N} L={L}
MPinv out n_nand vdd vdd    pfet_simple W={W_P} L={L}

* Charge sur la vraie sortie
CL out 0 10f

* ============================================
* Signal d'entrée
* ============================================
VIN in 0 PWL(
+ 0ns      0
+ 1ns      0
+ 1.02ns  {VDD_VAL}
+ 3ns     {VDD_VAL}
+ 3.02ns  0
+ 5ns     0
+ )

* ============================================
* Analyse transitoire et MESURES
* ============================================
.tran 0.01n 5.5n

* On mesure entre "in" et "out" (la sortie de l'inverseur)
* Note: Pour une porte AND, quand l'entrée monte, la sortie monte !
.measure tran tpLH TRIG v(in) VAL={VDD_VAL/2} RISE=1 TARG v(out) VAL={VDD_VAL/2} RISE=1
.measure tran tpHL TRIG v(in) VAL={VDD_VAL/2} FALL=1 TARG v(out) VAL={VDD_VAL/2} FALL=1
.measure tran tp PARAM='(tpLH + tpHL) / 2'

* Puissance
.measure tran I_stat FIND I(VVDD) AT=0.5n
.measure tran p_static PARAM='abs(I_stat)*VDD_VAL'
.measure tran Q_total INTEG I(VVDD) FROM=1n TO=5n
.measure tran E_total PARAM='abs(Q_total)*VDD_VAL'
.measure tran p_total PARAM='E_total/4n'
.measure tran p_dynamic PARAM='abs(p_total - p_static)'

.control
    run
    print tp p_static p_dynamic
    quit
.endc
.end
